`define ADDR_WIDTH 8
`define DATA_WIDTH 8
`define MEM_DEPTH 256
`define PSTRB_WIDTH 32
