`define ADDR_WIDTH 8
`define DATA_WIDTH 16
`define MEM_DEPTH 256
